library verilog;
use verilog.vl_types.all;
entity right_shift_8bit_vlg_vec_tst is
end right_shift_8bit_vlg_vec_tst;
