library verilog;
use verilog.vl_types.all;
entity booth_multiplier_8bit_vlg_vec_tst is
end booth_multiplier_8bit_vlg_vec_tst;
