library verilog;
use verilog.vl_types.all;
entity register_8bit_vlg_vec_tst is
end register_8bit_vlg_vec_tst;
