library verilog;
use verilog.vl_types.all;
entity register_vlg_check_tst is
    port(
        reg_output      : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end register_vlg_check_tst;
