library verilog;
use verilog.vl_types.all;
entity ripple_counter_4bit_vlg_vec_tst is
end ripple_counter_4bit_vlg_vec_tst;
