library verilog;
use verilog.vl_types.all;
entity mux4to1_16bit_vlg_vec_tst is
end mux4to1_16bit_vlg_vec_tst;
