library verilog;
use verilog.vl_types.all;
entity Sub_8bit_vlg_vec_tst is
end Sub_8bit_vlg_vec_tst;
