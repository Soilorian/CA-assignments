library verilog;
use verilog.vl_types.all;
entity gather_vlg_vec_tst is
end gather_vlg_vec_tst;
