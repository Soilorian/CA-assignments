library verilog;
use verilog.vl_types.all;
entity myALU_vlg_vec_tst is
end myALU_vlg_vec_tst;
