library verilog;
use verilog.vl_types.all;
entity register_2bit_vlg_vec_tst is
end register_2bit_vlg_vec_tst;
